// module operation
// p(x) = x^163 + x^80 + x^47 + x^9 + 1
module modulo(input [324:0]a,
              output [162:0]out);

    // maximum delay = 7 XOR gates
    assign out[7:0]     = a[7:0] ^ a[170:163] ^ a[324:317] ^ a[286:279] ^ a[253:246];
    assign out[8]       = a[8] ^ a[171] ^ a[287] ^ a[254];
    assign out[16:9]    = a[16:9] ^ a[179:172] ^ a[170:163] ^ a[324:317] ^ a[295:288] ^ a[286:279] ^ a[262:255] ^ a[253:246];
    assign out[45:17]   = a[45:17] ^ a[208:180] ^ a[199:171] ^ a[324:296] ^ a[315:287] ^ a[291:263] ^ a[282:254];
    assign out[46]      = a[46] ^ a[209] ^ a[200] ^ a[316] ^ a[292] ^ a[283];
    assign out[78:47]   = a[78:47] ^ a[241:210] ^ a[232:201] ^ a[194:163] ^ a[310:279] ^ a[324:293] ^ a[315:284] ^ a[277:246];
    assign out[79]      = a[79] ^ a[242] ^ a[233] ^ a[195] ^ a[311] ^ a[316] ^ a[278];
    assign out[92:80]   = a[92:80] ^ a[255:243] ^ a[246:234] ^ a[208:196] ^ a[175:163] ^ a[324:312] ^ a[258:246];
    assign out[158:93]  = a[158:93] ^ a[321:256] ^ a[312:247] ^ a[274:209] ^ a[241:176] ^ a[324:259]; 
    assign out[161:159] = a[161:159] ^ a[324:322] ^ a[315:313] ^ a[277:275] ^ a[244:242];
    assign out[162]     = a[162] ^ a[316] ^ a[278] ^ a[245];

endmodule