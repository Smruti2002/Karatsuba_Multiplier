module karatsuba_11x11(input [10:0]a,
                       input [10:0]b,
                       output [20:0]c);
    // normal multiplication
    
    assign c[0]  = a[0]&b[0];
    assign c[1]  = (a[0]&b[1]) ^ (a[1]&b[0]);
    assign c[2]  = (a[0]&b[2]) ^ (a[1]&b[1]) ^ (a[2]&b[0]);
    assign c[3]  = (a[0]&b[3]) ^ (a[1]&b[2]) ^ (a[2]&b[1]) ^ (a[3]&b[0]);
    assign c[4]  = (a[0]&b[4]) ^ (a[1]&b[3]) ^ (a[2]&b[2]) ^ (a[3]&b[1]) ^ (a[4]&b[0]);
    assign c[5]  = (a[0]&b[5]) ^ (a[1]&b[4]) ^ (a[2]&b[3]) ^ (a[3]&b[2]) ^ (a[4]&b[1]) ^ (a[5]&b[0]);
    assign c[6]  = (a[0]&b[6]) ^ (a[1]&b[5]) ^ (a[2]&b[4]) ^ (a[3]&b[3]) ^ (a[4]&b[2]) ^ (a[5]&b[1]) ^ (a[6]&b[0]);
    assign c[7]  = (a[0]&b[7]) ^ (a[1]&b[6]) ^ (a[2]&b[5]) ^ (a[3]&b[4]) ^ (a[4]&b[3]) ^ (a[5]&b[2]) ^ (a[6]&b[1]) ^ (a[7]&b[0]);
    assign c[8]  = (a[0]&b[8]) ^ (a[1]&b[7]) ^ (a[2]&b[6]) ^ (a[3]&b[5]) ^ (a[4]&b[4]) ^ (a[5]&b[3]) ^ (a[6]&b[2]) ^ (a[7]&b[1]) ^ (a[8]&b[0]);
    assign c[9]  = (a[0]&b[9]) ^ (a[1]&b[8]) ^ (a[2]&b[7]) ^ (a[3]&b[6]) ^ (a[4]&b[5]) ^ (a[5]&b[4]) ^ (a[6]&b[3]) ^ (a[7]&b[2]) ^ (a[8]&b[1]) ^ (a[9]&b[0]);
    assign c[10] = (a[0]&b[10]) ^ (a[1]&b[9]) ^ (a[2]&b[8]) ^ (a[3]&b[7]) ^ (a[4]&b[6]) ^ (a[5]&b[5]) ^ (a[6]&b[4]) ^ (a[7]&b[3]) ^ (a[8]&b[2]) ^ (a[9]&b[1]) ^ (a[10]&b[0]);
    assign c[11] = (a[1]&b[10]) ^ (a[2]&b[9]) ^ (a[3]&b[8]) ^ (a[4]&b[7]) ^ (a[5]&b[6]) ^ (a[6]&b[5]) ^ (a[7]&b[4]) ^ (a[8]&b[3]) ^ (a[9]&b[2]) ^ (a[10]&b[1]);
    assign c[12] = (a[2]&b[10]) ^ (a[3]&b[9]) ^ (a[4]&b[8]) ^ (a[5]&b[7]) ^ (a[6]&b[6]) ^ (a[7]&b[5]) ^ (a[8]&b[4]) ^ (a[9]&b[3]) ^ (a[10]&b[2]);
    assign c[13] = (a[3]&b[10]) ^ (a[4]&b[9]) ^ (a[5]&b[8]) ^ (a[6]&b[7]) ^ (a[7]&b[6]) ^ (a[8]&b[5]) ^ (a[9]&b[4]) ^ (a[10]&b[3]);
    assign c[14] = (a[4]&b[10]) ^ (a[5]&b[9]) ^ (a[6]&b[8]) ^ (a[7]&b[7]) ^ (a[8]&b[6]) ^ (a[9]&b[5]) ^ (a[10]&b[4]);
    assign c[15] = (a[5]&b[10]) ^ (a[6]&b[9]) ^ (a[7]&b[8]) ^ (a[8]&b[7]) ^ (a[9]&b[6]) ^ (a[10]&b[5]);
    assign c[16] = (a[6]&b[10]) ^ (a[7]&b[9]) ^ (a[8]&b[8]) ^ (a[9]&b[7]) ^ (a[10]&b[6]);
    assign c[17] = (a[7]&b[10]) ^ (a[8]&b[9]) ^ (a[9]&b[8]) ^ (a[10]&b[7]);
    assign c[18] = (a[8]&b[10]) ^ (a[9]&b[9]) ^ (a[10]&b[8]);
    assign c[19] = (a[9]&b[10]) ^ (a[10]&b[9]);
    assign c[20] = (a[10]&b[10]);

endmodule