`include "karatsuba_163.v"

module tb;

    reg [162:0]a;
    reg [162:0]b;
    wire [162:0]c;

    karatsuba_163x163 k(a,b,c);

    initial begin

        $monitor("c = %h\n",c);

        // test cases given in assignment
        a = 163'h8000000000000000000000000000000000000001;
        b = 163'h8000000000000000000000000000000000000001;
        #10;
        a = 163'h810000000000000000000000000000000000001;
        b = 163'h820000000000000000000000000000000000001;
        #10;
        a = 163'h7ffffffffffffffffffffffffffffffffffffffff;
        b = 163'h7ffffffffffffffffffffffffffffffffffffffff;
        #10;

        // x * (x^162) = 1 + x^9 + x^47 + x^80
        a = 163'h2;
        b = 163'h40000000000000000000000000000000000000000;
        #10;

        // x^162 * x^84 = 1 + x^9 + x^47 + x^80 + x^83 + x^92 + x^130
        a = 163'h40000000000000000000000000000000000000000;
        b = 163'h1000000000000000000000;
        #10;

        // x^162 * x^117 = 1 + x^9 + x^33 + x^42 + x^47 + x^113 + x^116 + x^125
        a = 163'h40000000000000000000000000000000000000000;
        b = 163'h200000000000000000000000000000;
        #10;
    end

endmodule 